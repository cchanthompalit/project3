library ieee;
use ieee.std_logic_1164.all;

package project_pkg is
    component Max10_adc is
        port (
            pll_clk:    in std_logic;
            chsel:      in natural range 0 to 2**5 - 1;
            soc:        in std_logic;
            tsen:       in std_logic;
            dout:       out natural range 0 to 2**12 - 1;
            eoc:        out std_logic;
            clk_dft:    out std_logic
        );
    end component Max10_adc;

    component synchronizer is
        generic (
            data_width: natural := 4
        );
        port (
            clk_a: in std_logic;
				clk_b: in std_logic;
            rst: in std_logic;
            data_in: in std_logic_vector(data_width - 1 downto 0);
            data_out: out std_logic_vector(data_width - 1 downto 0)
        );
    end component synchronizer;

    component bin_to_gray is
        generic (
            input_width: positive := 16
        );
        port (
            bin_in: in std_logic_vector(input_width - 1 downto 0);
            gray_out: out std_logic_vector(input_width - 1 downto 0)
        );
    end component bin_to_gray;

    component gray_to_bin is
        generic (
            input_width: positive := 16
        );
        port (
            gray_in: in std_logic_vector(input_width - 1 downto 0);
            bin_out: out std_logic_vector(input_width - 1 downto 0)
        );
    end component gray_to_bin;

    component true_dual_port_ram_dual_clock is
        generic (
            DATA_WIDTH : natural := 8;
            ADDR_WIDTH : natural := 6
        );
        port (
            clk_a: in std_logic; -- Single clock
				clk_b: in std_logic; -- Single clock
            addr_a: in natural range 0 to 2**ADDR_WIDTH - 1;
            addr_b: in natural range 0 to 2**ADDR_WIDTH - 1;
            data_a: in std_logic_vector((DATA_WIDTH-1) downto 0);
            data_b: in std_logic_vector((DATA_WIDTH-1) downto 0);
            we_a: in std_logic := '1';
            we_b: in std_logic := '1';
            q_a: out std_logic_vector((DATA_WIDTH -1) downto 0);
            q_b: out std_logic_vector((DATA_WIDTH -1) downto 0)
        );
    end component true_dual_port_ram_dual_clock;

    component adc_producer is
        generic (
            ADDR_WIDTH : natural := 6
        );
        port (
            clock: in std_logic; -- Single clock
            reset: in std_logic;
            tail_ptr: in natural range 0 to 2**ADDR_WIDTH - 1;
            eoc: in std_logic;
            soc: out std_logic;
            buffer_write: out std_logic;
            head_ptr: buffer natural range 0 to 2**ADDR_WIDTH - 1
        );
    end component adc_producer;

    component adc_control is
        generic (
            ADDR_WIDTH : natural := 6
        );
        port (
            clock: in std_logic; -- Single clock
            reset: in std_logic;
            head_ptr: in natural range 0 to 2**ADDR_WIDTH - 1;
            tail_ptr: buffer natural range 0 to 2**ADDR_WIDTH - 1
        );
    end component adc_control;

    component pll is
        port (
            inclk0: in STD_LOGIC := '0';
            c0: OUT STD_LOGIC 
        );
    end component pll;

end package project_pkg;
